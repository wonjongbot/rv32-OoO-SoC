`define PROJECT_ROOT "/home/wonjongbot/rv32-OoO-SoC/"
